`define data_width 8
`define addr_width 9
